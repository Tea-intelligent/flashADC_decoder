`timescale 1ns/1ps
module tb();
integer     fd; 
reg [254:0]data_I;
wire [7:0]data_O;


initial begin 
fd = $fopen("output.txt","w");
data_I=255'd0;
#10
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");
data_I=255'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
#10;
$fwrite(fd, data_O);
$fwrite(fd, "\n");





#2000 $finish;

end
final f_instance(.O(data_O),.In(data_I));

endmodule
